`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2020/01/12 21:49:01
// Design Name: 
// Module Name: pd_sim
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module pd_sim(

    );
    
//    reg [7:0] clk;
//    reg [255:0] data;
//    wire sig;
//    wire clk_out;
//    phase_detector #(8)
//    pd(clk,sig,clk_out);
//    initial clk<=8'hf0;
//    initial data<=256'h136F855C63C94DC3F1237E253FB42F8ADB7B3011C0AB13F224478C6A0F409879;
//    always #2 clk<={clk[6:0],clk[7]};
//    initial #1 forever #8 repeat(16) #16 data<={data[0],data[255:1]};
//    assign sig=data[0];
//    initial #4096 $finish;
endmodule
